class driver extends uvm_driver;
	function new(string name="driver", uvm_component parent);
	super.new(name,parent);
endfunction
endclass
