class monitor extends uvm_monitor;
endclass
