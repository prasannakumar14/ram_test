class monitor extends uvm_monitor;
	function new(string name="monitor", uvm_component parent);
		super.new(name,parent);
	endfunction
endclass
